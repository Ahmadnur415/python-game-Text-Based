��M	      �game_rpg.game��Game���)��}�(�player��game_rpg.player��Player���)��}�(�strength�K�magic�K�archery�K�constitution�K
�will�K�
perception�K�	growth_hp�KZ�	growth_mp�Kx�luck�KZ�defense�K�evasion�K�
resistance�K1�armor_penetration�K�_max_health�K}�	_max_mana�K�_max_stamina�K�_health�K��_mana�K�_stamina�K�_Entity__name��Ahmad��_Entity__namespace��player��_Entity__class��mage��level�K�	equipment�}�(�	main_hand��game_rpg.items.items��Items���)��}�(�name��magic wood staff��quality�K �	typeItems��weapons��identify��staff:m_staff��	attribute�h(�
EQUIPPABLE���)��}�(�use���location�]��	main_hand�a�user�]��mage�a�styleAttack��game_rpg.attack��_attackstyle���)��}��damage_stats��magic�sb�attack�]�hA�Attack���)��}�(h-�magic:magicbolt��displayName��
magic bolt��
typeAttack��magic��base_damage�]�(KKe�description_of_being_used��fire an magic bolt at��cost_mp�K�cost_st�K �effect�]��
multiplier�]�(hA�
Multiplier���)��}�(�modifier�G?ə������stats��
self.magic�ubh^)��}�(haG?�      hb�self.magic_damage�ubeuba�
classItems��staff��damage�hThKhK hK hK ub�amount�K�price�}�(�value�Kd�type��silver��max_discount�K u�	sub_stats�}�(�magic�K�will�K�
perception�J����u�in_shop��ub�off_hand�N�two_hand�N�head�N�body�h*)��}�(h-�Saint's Robe�h/K h0�armor�h2�armor:saints_r�h4h6)��}�(h9�h:]��body�ah=�all�h@NhH]�hg�armor�hiK hK hK hKhK ubhjKhk}�(�value�M��type��silver��max_discount�Kuhq}�hv�ub�shoes�h*)��}�(h-�Gardener Shoes�h/K h0�armor�h2�footgear:gardener_shoes�h4h6)��}�(h9�h:]��shoes�ah=]��all�ah@NhH]�hg�footgear�hiK hK hKhK
hK ubhjKhk}�(�value�Kd�type��silver��max_discount�K uhq}��health�Kdshv�ubu�	inventory�]�(h+h�h{h*)��}�(h-�Blue Potion�h/Kh0�potion�h2�potion:blue_potion�h4h(�
CONSUMABLE���)��}�(hY]��type_��restore�hb}��mana�}�(�value�K�modiefer��max_mana�usubhjKhk}�(h�K#�type��silver��max_discount�K uhq}�ubehH]�(hK)��}�(h-�basic_attack:03�hO�Basic Attack�hQ�physical�hS]�(KK	ehU�attack�hWK hXK hY]�h[]�(h^)��}�(haG?�      hb�
self.level�ubh^)��}�(haG?�333333hb�self.physical_damage�ubh^)��}�(haG?ٙ�����hb�
self.magic�ubeubhLe�type_attack��magic��style_attack��magic��silver�JH� �gold�J�B �exp�K<�point_level�K�setting�}�ubh�}�(�	auto_gave���input_prompt��>>> ��lang��en_US��
difficulty�K�savename��Ahmad.sv�uub.
���      �game_rpg.game��Game���)��}�(�player��game_rpg.player��Player���)��}�(�strength�K#�magic�K�archery�K#�constitution�K�will�K�
perception�K�	growth_hp�K_�	growth_mp�Ki�luck�Kx�defense�MM�evasion�K�
resistance�K�armor_penetration�Km�_max_health�K�_max_stamina�KK�	_max_mana�K
�_health�KQ�_mana�K"�_stamina�K'�_Entity__name��body��_Entity__namespace��player��_Entity__class��archer��level�K�	equipment�}�(�	main_hand�N�off_hand�N�two_hand��game_rpg.items.items��Items���)��}�(�name��Bow Of Storm��quality�K�	typeItems��weapons��identify��bow:bow_of_storm��	attribute�h*�
EQUIPPABLE���)��}�(�use���location�]��two_hand�a�user�]��archer�a�styleAttack��game_rpg.attack��_attackstyle���)��}��damage_stats��archery�sb�attack�]�(hC�Attack���)��}�(h/�ranged:shoot��displayName��shoot��
typeAttack��physical��base_damage�]�(KKe�description_of_being_used��Shoot at��cost_mp�K �cost_st�K�effect�]��
multiplier�]�(hC�
Multiplier���)��}�(�modifier�G?ə������stats��self.magic_damage�ubh`)��}�(hcG?�ffffffhd�self.damage�ubeubhM)��}�(h/�ranged:one_shoot�hQ�	one shoot�hS�physical�hU]�(KK
ehWhXhYK hZK2h[]�h]]�(h`)��}�(hcG?�������hd�
self.level�ubh`)��}�(hcG?�      hd�enemy.archery�ubh`)��}�(hcG?�      hd�self.damage�ubeube�
classItems��bow��damage�hnhKdhK hK hK ub�amount�K�price�}�(�value�M��type��gold��max_discount�K u�	sub_stats�}�(�stamina�K2�critical_hit�Kdu�in_shop��ub�head�h,)��}�(h/�	King helm�h1Kh2�armor�h4�helmet:king_helm�h6h8)��}�(h;�h<]��head�ah?�all�hBNhJ]�hz�helmet�h|K hK hKhKhK ubh}Kh~}�(�value�K�type��gold��max_discount�Kuh�}�(�constitution�K�strength�K�will�Kuh��ub�body�h,)��}�(h/�Legendaty Armor�h1Kh2�armor�h4�armor:l_armor�h6h8)��}�(h;�h<]��body�ah?�all�hBNhJ]�hz�armor�h|K hK hK�hK
hK ubh}Kh~}�(�value�Kc�type��gold��max_discount�Kuh�}�(�constitution�K
�will�K
�
perception�K
uh��ub�shoes�h,)��}�(h/�Battle Boots�h1Kh2�armor�h4�footgear:battle_boots�h6h8)��}�(h;�h<]��shoes�ah?]��all�ahBNhJ]�hz�footgear�h|K hK hK6hK hK ubh}Kh~}�(�value�Kd�type��gold��max_discount�Kuh�}�(�strength�K�magic�K�archery�Kuh��ubu�	inventory�]�(h,)��}�(h/�
Wooden Bow�h1K h2h3h4�
bow:wood_b�h6h8)��}�(h;�h<h=h?h@hBhFhJ]�hM)��}�(h/hPhQhRhShThUhVhWhXhYK hZKh[]�h]]�(h`)��}�(hcG?ə�����hdheubh`)��}�(hcG?�ffffffhdhhubeubahzh{h|]�(KK
ehKhK hK hK ubh}Kh~}�(h�Kdh��silver�h�K uh�}�(�archery�K�critical_change�Kuh��ubh,)��}�(h/�Saint's Robe�h1K h2h�h4�armor:saints_r�h6h8)��}�(h;�h<h�h?h�hBNhJ]�hzh�h|K hK hK hKhK ubh}Kh~}�(h�M�h��silver�h�Kuh�}�h��ubh,)��}�(h/�Recover Potion�h1K h2�potion�h4�potion:recover_potion�h6h*�
CONSUMABLE���)��}�(h[]��type_��restore�hd}�(�health�K
�mana�K2�stamina�Kuubh}Kh~}�(�value�K��type��silver��max_discount�Kuh�}�ubh�h�h-h�h,)��}�(h/�Assassin Mask�h1K h2h�h4�helmet:assassin_mask�h6h8)��}�(h;�h<h�h?h�hBNhJ]�hzh�h|K hK hK hK hK ubh}Kh~}�(h�M�h��silver�h�K uh�}�(�critical_change�K�critical_hit�K
uh��ubehJ]�(hM)��}�(h/�basic_attack:02�hQ�Basic Attack�hS�physical�hU]�(KK
ehW�attack�hYK hZK h[]�h]]�(h`)��}�(hcG?�      hd�
self.level�ubh`)��}�(hcG?�333333hd�self.physical_damage�ubh`)��}�(hcG?ٙ�����hd�self.archery�ubeubhNhie�type_attack��physical��style_attack��archery��silver�Jr� �gold�J�? �exp�M'�point_level�K�setting�}�ubj*  }�(�	auto_gave���input_prompt��>>> ��lang��en_US��
difficulty�K�savename��body.sv�uub.